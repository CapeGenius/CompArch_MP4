module mux3 #(parameter WIDTH=32)
    (
        // Three data lines
        input logic [WIDTH - 1: 0] d0,
        input logic [WIDTH - 1: 0] d1,
        input logic [WIDTH - 1: 0] d2,
        
        // Select channel
        input logic [1:0] s,

        // Output selected data
        output logic [WIDTH - 1: 0] y
    );

    assign y = s[1] ? d2 : (s[0] ? d1 : d0);
endmodule
